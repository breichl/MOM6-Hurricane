.datasets/OM4_0p25_JR55/INPUTS/hycom1_75.cdl