.datasets/OM4_0p25_JR55/INPUTS/Oman_RedSea.cdl