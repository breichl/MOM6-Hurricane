.datasets/OM4_0p25_JR55/INPUTS/Faroe_GS_edits.cdl