.datasets/OM4_0p25_JR55/INPUTS/analysis_vgrid_lev35.v1.cdl