.datasets/OM4_0p25_JR55/INPUTS/Wyville_Thompson_edits.cdl