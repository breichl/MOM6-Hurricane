.datasets/OM4_0p25_JR55/INPUTS/Caribbean_edits.cdl