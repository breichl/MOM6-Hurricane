.datasets/OM4_0p25_JR55/INPUTS/vgrid_75_2m_575m.cdl